`include "ram_tx.sv"
`include "ram_gtr.sv"
`include "ram_drv.sv"
`include "ram_mon.sv"
`include "ram_refer.sv"
`include "ram_sb.sv"
`include "ram_env.sv"
`include "ram_test.sv"
