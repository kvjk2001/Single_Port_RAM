`include "../rtl/ram_design.v"
`include "ram_interface.sv"
`include "ram_sequence_item.sv"
`include "ram_sequence.sv"
`include "ram_sequencer.sv"
`include "ram_driver.sv"
`include "ram_in_monitor.sv"
`include "ram_active_agent.sv"
`include "ram_out_monitor.sv"
`include "ram_passive_agent.sv"
`include "ram_coverage.sv"
`include "ram_reference.sv"
`include "ram_scoreboard.sv"
`include "ram_environment.sv"
`include "ram_test.sv"
