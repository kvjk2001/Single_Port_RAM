`timescale 1ns/100ps

`define DATA_WIDTH 8
`define DATA_DEPTH 32
`define num_transactions 10
`define ADDR_WIDTH 5
