`include "../rtl/ram_design.v"
`include "intf.sv"
`include "sequence_item.sv"
`include "sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "in_monitor.sv"
`include "active_agent.sv"
`include "out_monitor.sv"
`include "passive_agent.sv"
`include "coverage.sv"
`include "reference.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"
