`define width 8
`define depth 256

`define no_of_seq 1
