`define no_of_seq 1
